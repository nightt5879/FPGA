`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: lab1
//////////////////////////////////////////////////////////////////////////////////

module lab1(
    input [3:0] swt,  // 修改为4个输入开关
    output [3:0] led  // 修改为4个输出 LED
    );

    // 逻辑更改成直接每个LED对应每一个按键
    // 需要注意的是按下按键是低电平，LED也是低电平亮灯，具体原因可以自行查阅数据手册
    assign led[0] = swt[0];                
    assign led[1] = swt[1];       
    assign led[2] = swt[2];        
    assign led[3] = swt[3];        

endmodule
